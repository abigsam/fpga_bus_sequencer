`ifndef __BUS_SEQUENCER_BASIC_TEST_SV
`define __BUS_SEQUENCER_BASIC_TEST_SV

class bus_sequencer_basic_test extends uvm_test;

    //**************************************************************************
    //declaring component utils for the basic test-case 
    //**************************************************************************
    `uvm_component_utils(bus_sequencer_basic_test)


    //**************************************************************************
    // Method name : new
    // Decription: Constructor 
    //**************************************************************************
    function new(string name = "bus_sequencer_basic_test",uvm_component parent=null);
        super.new(name,parent);
    endfunction : new

    //**************************************************************************
    // Method name : build_phase
    // Decription: Construct the components and objects
    //**************************************************************************
    virtual function void build_phase(uvm_phase phase);
        super.build_phase(phase);

        env = bus_sequencer_environment::type_id::create("env", this);
        seq = bus_sequencer_basic_seq::type_id::create("seq");
    endfunction : build_phase

    //**************************************************************************
    // Method name : run_phase
    // Decription: Trigger the sequences to run
    //**************************************************************************
    task run_phase(uvm_phase phase);
        phase.raise_objection(this);
        seq.start(env.bus_sequencer_agnt.sequencer);
        phase.drop_objection(this);
    endtask : run_phase

endclass : bus_sequencer_basic_test

`endif //__BUS_SEQUENCER_BASIC_TEST_SV