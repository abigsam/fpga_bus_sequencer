`ifndef __BUS_SEQUENCER_TB_TOP_SV
`define __BUS_SEQUENCER_TB_TOP_SV

`include "uvm_macros.svh"
`include "bus_sequencer_interface.sv"

import uvm_pkg::*;

module bus_sequencer_tb_top;

    import bus_sequencer_test_list::*;


    //**************************************************************************

    //**************************************************************************



endmodule

`endif //__BUS_SEQUENCER_TB_TOP